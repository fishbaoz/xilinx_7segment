//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    19:38:17 07/21/2008
// Design Name:
// Module Name:    ila_4kx32
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module ila_4kx32  (
    input [35:0] control,
    input clk,
    input [31:0] data,
    input [31:0] trig0
    );
endmodule

