//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    19:37:46 07/21/2008
// Design Name:
// Module Name:    icon
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

/******************************************************************************
 ***       the ICON hardmacro module onion skin                             ***
 ******************************************************************************/
module icon (
    input tdo_in,
    output tdi_out,
    output reset_out,
    output shift_out,
    output update_out,
    output sel_out,
    output drck_out,
    output [35:0] control0
    );
endmodule

